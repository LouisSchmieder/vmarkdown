module main

import parser

fn main() {
	mut parser := parser.new_parser('# Hello there')
}